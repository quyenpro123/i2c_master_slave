program testcase();

endprogram