`ifndef SCB
`define SCB
class scoreboard;
    logic [7:0] slave_addr;
    logic [7:0] data;
endclass
`endif