module top_tb (
    ports
);
    
endmodule