class assertion;
    
endclass //className