module i2c_fifo_block(
    
);


endmodule