////////////////////////////////////////////////
////s~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~s////
////s           www.testbench.in           s////
////s                                      s////
////s        SystemVerilog Tutorial        s////
////s                                      s////
////s           gopi@testbench.in          s////
////s~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~s////
////////////////////////////////////////////////
`ifndef INTF
`define INTF


interface intf_cnt(input logic pclk, input logic i2c_core_clock);
    //input dut
    logic preset;
    logic [7:0] paddr;
    logic pwrite;
    logic psel;
    logic penable;
    logic [7:0] pwdata;
    //output dut
    wire sda_io;
    wire scl_io;
    logic [7:0] prdata_o;
    logic pready_o;
    logic stop;
    logic start;
endinterface
`endif
