class monitor;

endclass