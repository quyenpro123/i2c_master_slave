`ifndef MOR
`define MOR 
class monitor;

endclass
`endif