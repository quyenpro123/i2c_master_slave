class environment;

endclass