class transactor;
    rand logic [7:0]    pwdata;
    rand logic [7:0]    paddr;
    rand logic          pwrite;
    rand logic          psel;
    rand logic          penable;
endclass //transactor